class env_config extends uvm_object;

function new(string name = "env_config");
    super.new(name);
endfunction

bit has_scb = 1;

endclass
