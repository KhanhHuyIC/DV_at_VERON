module ha_1b (
  input
