`timescale 1ns/1ps

//====================== Interface ======================//
interface fifo_if #(parameter DATA_WIDTH = 8) ();
    logic clk;                             // Clock signal
    logic rst_n;                           // Active low reset signal
    logic wr, rd, clear;                   // Write, read, and clear signals
    logic [DATA_WIDTH-1:0] data_in;        // Input data to be written
    logic data_out_valid;                  // Valid output data signal
    logic [DATA_WIDTH-1:0] data_out;       // Output data read from FIFO
    logic empty, full;                     // FIFO empty and full flags
endinterface


//=================== Transaction =======================//
class FIFO_transaction #(parameter DATA_WIDTH = 8);
    // Data members
    bit wr;                            // Write signal
    bit rd;                            // Read signal
    bit [DATA_WIDTH-1:0] data;         // Data associated with the transaction

    // Constructor
    function new(input bit wr, input bit rd, input [DATA_WIDTH-1:0] data);
        this.wr = wr;
        this.rd = rd;
        this.data = data;
    endfunction

    // Print Method for debugging
    function void print();
        $display("Write: %b, Read: %b, Data: %h", wr, rd, data);
    endfunction
endclass


//==================== Generator ========================//
class FIFO_generator #(parameter DATA_WIDTH = 8);
    mailbox #(FIFO_transaction #(DATA_WIDTH)) gen2drv;

    virtual fifo_if #(DATA_WIDTH) vif;

    function new(mailbox #(FIFO_transaction #(DATA_WIDTH)) gen2drv, virtual fifo_if #(DATA_WIDTH) vif);
        this.gen2drv = gen2drv;
        this.vif = vif;
    endfunction

    task run();
    FIFO_transaction #(DATA_WIDTH) tr;

    // --- Step 1: Write a few samples
    for (int i = 0; i < 5; i++) begin
        tr = new(1, 0, $urandom_range(0, 255));
        gen2drv.put(tr);
        tr.print();
        #20;
    end

    // --- Step 2: Idle for a few cycles
    for (int i = 0; i < 3; i++) begin
        tr = new(0, 0, 8'h00);
        gen2drv.put(tr);
        #20;
    end

    // --- Step 3: Read a few samples
    for (int i = 0; i < 3; i++) begin
        tr = new(0, 1, 8'h00);
        gen2drv.put(tr);
        tr.print();
        #20;
    end

    // --- Step 4: Write continuously until FIFO is full
    while (vif.full !== 1) begin
        tr = new(1, 0, $urandom_range(0, 255));
        gen2drv.put(tr);
        tr.print();
        #20;
    end
    $display("[GEN] FIFO FULL detected, stop writing");

    // --- Step 5: Read a few samples from FIFO
    for (int i = 0; i < 4; i++) begin
        tr = new(0, 1, 8'h00);
        gen2drv.put(tr);
        tr.print();
        #20;
    end

    // --- Step 6: Idle again for a few cycles
    for (int i = 0; i < 3; i++) begin
        tr = new(0, 0, 8'h00);
        gen2drv.put(tr);
        #20;
    end

    // --- Step 7: Read continuously until FIFO is empty
    while (vif.empty !== 1) begin
        tr = new(0, 1, 8'h00);
        gen2drv.put(tr);
        tr.print();
        #20;
    end
    $display("[GEN] FIFO EMPTY detected, stop reading");
    endtask

endclass


//====================== Driver =========================//
class FIFO_driver #(parameter DATA_WIDTH = 8);
    virtual fifo_if #(DATA_WIDTH) vif;                 // Virtual interface to connect with the DUT
    mailbox #(FIFO_transaction #(DATA_WIDTH)) gen2drv; // Mailbox to receive transactions from the generator

    // Constructor to initialize the driver
    function new(virtual fifo_if #(DATA_WIDTH) vif, mailbox #(FIFO_transaction #(DATA_WIDTH)) gen2drv);
        this.vif = vif;              // Connect virtual interface to the DUT
        this.gen2drv = gen2drv;      // Connect the mailbox to receive transactions
    endfunction

    // Task to drive signals based on the received transaction
    task run();
        FIFO_transaction #(DATA_WIDTH) tr;  // Transaction object to store incoming data
        forever begin
            gen2drv.get(tr);  // Get a transaction from the mailbox (generated by the generator)

            @(posedge vif.clk);  // Wait for the rising edge of the clock
            vif.wr      <= tr.wr;  // Drive the write signal
            vif.rd      <= tr.rd;  // Drive the read signal
            vif.data_in <= tr.data;  // Drive the data input signal

            @(posedge vif.clk);  // Wait for another rising clock edge
            vif.wr <= 0;  // Reset write signal
            vif.rd <= 0;  // Reset read signal
            #10;  // Wait for a small delay before the next transaction
        end
    endtask

endclass



//===================== Monitor =========================//
class FIFO_monitor #(parameter DATA_WIDTH = 8);
    virtual fifo_if #(DATA_WIDTH) vif;                   // Virtual interface to observe DUT
    mailbox #(FIFO_transaction #(DATA_WIDTH)) mon2sb;    // Mailbox to send captured transactions to the scoreboard

    // Constructor to initialize the monitor
    function new(virtual fifo_if #(DATA_WIDTH) vif, mailbox #(FIFO_transaction #(DATA_WIDTH)) mon2sb);
        this.vif = vif;                // Connect virtual interface to the DUT for observation
        this.mon2sb = mon2sb;          // Connect mailbox to send captured data to the scoreboard
    endfunction

    // Task to monitor and capture outputs
    task run();
        FIFO_transaction #(DATA_WIDTH) tr;  // Transaction object to store captured data
        forever begin
            @(posedge vif.clk);  // Wait for the rising clock edge

            // Check if the write signal is active
            if (vif.wr) begin
                tr = new(1, 0, vif.data_in);  // Create a write transaction with the data_in value
                mon2sb.put(tr);  // Send the write transaction to the scoreboard
            end

            // Check if the data_out_valid signal is active
            if (vif.data_out_valid) begin
                tr = new(0, 1, vif.data_out);  // Create a read transaction with the data_out value
                mon2sb.put(tr);  // Send the read transaction to the scoreboard
            end
        end
    endtask

endclass

//==================== Scoreboard =======================//
class FIFO_scoreboard #(parameter DATA_WIDTH = 8);
    mailbox #(FIFO_transaction #(DATA_WIDTH)) mon2sb;
    bit [DATA_WIDTH-1:0] model[$];

    function new(mailbox #(FIFO_transaction #(DATA_WIDTH)) mon2sb);
        this.mon2sb = mon2sb;
    endfunction

    task run();
        FIFO_transaction #(DATA_WIDTH) tr;
        forever begin
            mon2sb.get(tr);
            if (tr.wr && !tr.rd) begin
                model.push_back(tr.data);
                $display("[SB] PUSH data=0x%0h", tr.data);
            end else if (!tr.wr && tr.rd) begin
                if (model.size() > 0) begin
                    bit [DATA_WIDTH-1:0] expected = model.pop_front();
                    $display("[SB] POP  expect=0x%0h", expected);
                end else begin
                    $display("[SB] ERROR: Read when FIFO empty");
                end
            end
        end
    endtask
endclass

//==================== Environment ======================//
class FIFO_env #(parameter DATA_WIDTH = 8);
    FIFO_generator #(DATA_WIDTH) gen;
    FIFO_driver    #(DATA_WIDTH) drv;
    FIFO_monitor   #(DATA_WIDTH) mon;
    FIFO_scoreboard #(DATA_WIDTH) sb;

    mailbox #(FIFO_transaction #(DATA_WIDTH)) gen2drv;
    mailbox #(FIFO_transaction #(DATA_WIDTH)) mon2sb;

    virtual fifo_if #(DATA_WIDTH) vif;

    function new(virtual fifo_if #(DATA_WIDTH) vif);
        this.vif = vif;
        gen2drv = new();
        mon2sb  = new();
        sb      = new(mon2sb);
        gen     = new(gen2drv, vif);
        drv     = new(vif, gen2drv);
        mon     = new(vif, mon2sb);
    endfunction

    task run();
        fork
            gen.run();
            drv.run();
            mon.run();
            sb.run();
        join_any
    endtask
endclass


//======================= Testbench Top ===========================//
module FIFO_8b_tb;
    fifo_if #(8) intf();

    // Clock generation
    initial begin
        intf.clk = 0;
        forever #5 intf.clk = ~intf.clk;
    end

    // Reset
    initial begin
        intf.wr = 0;
        intf.rd = 0;
        intf.data_in = 0;
        intf.rst_n = 0;
        intf.clear = 0;
        #12;
        intf.rst_n = 1;
    end

    //Test clear signal
    initial begin
    #525;
    $display("[TB] Trigger clear");
    intf.clear = 1;
    #20;
    intf.clear = 0;
    end

    // DUT instantiation
    FIFO_8b dut (
        .clk(intf.clk),
        .rst_n(intf.rst_n),
        .wr(intf.wr),
        .rd(intf.rd),
        .clear(intf.clear),
        .data_in(intf.data_in),
        .data_out_valid(intf.data_out_valid),
        .data_out(intf.data_out),
        .empty(intf.empty),
        .full(intf.full)
    );

    // Dump for waveform
    initial begin
        $dumpfile("fifo_8b_tb.vcd");
        $dumpvars(0, FIFO_8b_tb);
    end

    // Environment
    FIFO_env #(8) env;

    initial begin
        env = new(intf);
        $monitor($time, " wr=%b rd=%b data_in=%h data_out=%h valid=%b full=%b empty=%b",
                 intf.wr, intf.rd, intf.data_in, intf.data_out, intf.data_out_valid, intf.full, intf.empty);
        env.run();
        #2000;
        $finish;
    end

    //Simple assertion
    always @(posedge intf.clk) begin
    if (intf.rd && intf.empty)
        $error("ASSERT: Reading from empty FIFO!");

    if (intf.wr && intf.full)
        $error("ASSERT: Writing to full FIFO!");
    end

    //Simple Coverage
    integer wr_count = 0, rd_count = 0;

    always @(posedge intf.clk)
    if (intf.wr && !intf.full) wr_count++;

    always @(posedge intf.clk)
    if (intf.rd && intf.data_out_valid) rd_count++;

    final begin
        $display("[COV] Total write cycles: %0d", wr_count);
        $display("[COV] Total read cycles : %0d", rd_count);
    end

endmodule
